** Profile: "SCHEMATIC1-simprof"  [ C:\Users\dawnm\Desktop\Steilto\opamp-final\Operational Amplifier\opamp_final-pspicefiles\schematic1\simprof.sim ] 

** Creating circuit file "simprof.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
.LIB "../../../opamp_final-pspicefiles/opamp_final.lib" 
* From [PSPICE NETLIST] section of C:\Users\dawnm\AppData\Roaming\SPB_Data\cdssetup\OrCAD_PSpice\17.2.0\PSpice.ini file:
.lib "nomd.lib" 

*Analysis directives: 
.AC DEC 10 10 100meg
.OPTIONS ADVCONV
.PROBE64 V(*) I(*) W(*) D(*) NOISE(*) 
.INC "..\SCHEMATIC1.net" 


.END
